// Created by altera_lib_mf.pl from altera_mf.v

/*verilator lint_off CASEX*/
/*verilator lint_off COMBDLY*/
/*verilator lint_off INITIALDLY*/
/*verilator lint_off LITENDIAN*/
/*verilator lint_off MULTIDRIVEN*/
/*verilator lint_off UNOPTFLAT*/
/*verilator lint_off BLKANDNBLK*/
module    altstratixii_oct    (
    terminationenable,
    terminationclock,
    rdn,
    rup);

    parameter    lpm_type    =    "altstratixii_oct";


    input    terminationenable;
    input    terminationclock;
    input    rdn;
    input    rup;

endmodule //altstratixii_oct

